`timescale 1ns / 1ns // `timescale time_unit/time_precision


//code to display on hex0 and hex1
module hex7seg (input[3:0] c, output[0:6] led);

	assign led[0] = (~c[3]&~c[2]&~c[1]&c[0])|(~c[3]&c[2]&~c[1]&~c[0])|
						 (c[3]&~c[2]&c[1]&c[0])|(c[3]&c[2]&~c[1]&c[0]);
						  
	assign led[1] = (~c[3]&c[2]&~c[1]&c[0])|(~c[3]&c[2]&c[1]&~c[0])|
						 (c[3]&~c[2]&c[1]&c[0])|(c[3]&c[2]&~c[1]&~c[0])|
					    (c[3]&c[2]&c[1]&~c[0])|(c[3]&c[2]&c[1]&c[0]);
						  
	assign led[2] = (~c[3]&~c[2]&c[1]&~c[0])|(c[3]&c[2]&~c[1]&~c[0])|
						 (c[3]&c[2]&c[1]&~c[0])|(c[3]&c[2]&c[1]&c[0]);
	
	assign led[3] = (~c[3]&~c[2]&~c[1]&c[0])|(~c[3]&c[2]&~c[1]&~c[0])|
						 (~c[3]&c[2]&c[1]&c[0])|(c[3]&~c[2]&c[1]&~c[0])|
						 (c[3]&c[2]&c[1]&c[0]);
						  
	
	assign led[4] = (~c[3]&~c[2]&~c[1]&c[0])|(~c[3]&~c[2]&c[1]&c[0])|
						 (~c[3]&c[2]&~c[1]&~c[0])|(~c[3]&c[2]&~c[1]&c[0])|
						 (~c[3]&c[2]&c[1]&c[0])|(c[3]&~c[2]&~c[1]&c[0]);
						  
	
	assign led[5] = (~c[3]&~c[2]&~c[1]&c[0])|(~c[3]&~c[2]&c[1]&~c[0])|
						 (~c[3]&~c[2]&c[1]&c[0])|(~c[3]&c[2]&c[1]&c[0])|
						 (c[3]&c[2]&~c[1]&c[0]);
						  
	
	assign led[6] = (~c[3]&~c[2]&~c[1]&~c[0])|(~c[3]&~c[2]&~c[1]&c[0])|
						 (~c[3]&c[2]&c[1]&c[0])|(c[3]&c[2]&~c[1]&~c[0]);

endmodule
